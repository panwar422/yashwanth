module tb;
    initial 
    begin
        $display("hi");
    end
endmodule 